---------------------------------
--	State Machine for the LCD
--	driver
---------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY lcd IS 
	PORT(
		clk, rst : STD_LOGIC);
END lcd;

ARCHITECTURE behaviour OF lcd IS

BEGIN
	
END behaviour;
