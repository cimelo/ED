---------------------------------
--	State Machine for the LCD
--	driver
---------------------------------

ENTITY lcd IS 
	PORT(
		clk, rst : ST
	);
END lcd;

ARCHITECTURE behaviour OF lcd IS

BEGIN
	
END behaviour;
